module tb;
reg rst,clk;
wire sda;
reg scl;
reg lane;
reg [7:0] data_send_slave;
reg data_send_slave_enable;
wire [7:0] data_receive_slave;
wire data_receive_slave_enable;
wire error_slave;
assign sda=lane;

i2c_slave dut(
.rst(rst),
.clk(clk),
.scl(scl),.sda(sda),
.data_send_slave_enable(data_send_slave_enable),
.data_receive_slave_enable(data_receive_slave_enable),
.data_send_slave(data_send_slave),
.data_receive_slave(data_receive_slave),
.error_slave(error_slave)
);
initial begin
clk=1;
forever #5 clk=~clk;
#500;
$stop;
end
initial begin
	scl=1;
	#55;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#150;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
	scl=~scl;
	#10;
end
initial begin
	rst<=0;
	data_send_slave<=8'h00;
	data_send_slave_enable<=1'b0;
	lane<=1'b1;
	#20;
	rst<=1;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#20;
	lane=1'b0;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#20;
	lane=1'b1;
	#20;
	lane=1'b0;
	#20;
	lane=1'bz;
	#20;
	lane=1'b1;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#20;
	lane=1'b1;
	#20;
	lane=1'b1;
	#20;
	lane=1'b1;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#20;
	lane=1'bz;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#120;
	data_send_slave_enable=1'b1;
	data_send_slave=8'h93;
	lane=1'b0;
	#20;
	data_send_slave_enable=1'b0;
	data_send_slave=8'h00;
	lane=1'b1;
	#20;
	lane=1'b0;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#20;
	lane=1'b1;
	#20;
	lane=1'b1;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'bz;
	#20;
	lane=1'b0;
	#20;
	lane=1'b0;
	#20;
	lane=1'b1;
	#50;
	$stop;
end	
endmodule
